`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/06/2020 02:02:02 PM
// Design Name: 
// Module Name: fmul_pipelined
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module pipelined_fmul (a,b,rm,s,clk,clrn,e); // pipelined fp mul
    input [31:0] a, b; // fp a and b
    input [1:0] rm; // round mode
    input e; // enable
    input clk, clrn; // clock and reset
    output [31:0] s; // fp output
    
    wire m_sign;
    wire [9:0] m_exp10;
    wire m_is_nan;
    wire m_is_inf;
    wire [22:0] m_inf_nan_frac;
    wire [39:0] m_sum;
    wire [39:0] m_carry;
    wire [7:0] m_z8;
    // exe1: partial product stage (carry and sum generated by wallace tree)
    fmul_mul mul1 (a,b,m_sign,m_exp10,m_is_nan,m_is_inf,m_inf_nan_frac,m_sum,m_carry,m_z8);
    wire [1:0] a_rm;
    wire a_sign;
    wire [9:0] a_exp10;
    wire a_is_nan;
    wire a_is_inf;
    wire [22:0] a_inf_nan_frac;
    wire [39:0] a_sum;
    wire [39:0] a_carry;
    wire [7:0] a_z8;
    // pipeline register
    reg_mul_add reg_ma(rm,m_sign,m_exp10,m_is_nan,m_is_inf,m_inf_nan_frac,
                        m_sum,m_carry,m_z8,clk,clrn,e, a_rm,a_sign,a_exp10,
                        a_is_nan,a_is_inf,a_inf_nan_frac,a_sum,a_carry,a_z8);
    wire [47:8] a_z40;
    // exe2: addition stage (product by adding carry and sum)
    fmul_add mul2 (a_sum,a_carry,a_z40);
    wire [47:0] a_z48 = {a_z40,a_z8};
    wire [1:0] n_rm;
    wire n_sign;
    wire [9:0] n_exp10;
    wire n_is_nan;
    wire n_is_inf;
    wire [22:0] n_inf_nan_frac;
    wire [47:0] n_z48;
    // pipeline register
    reg_add_norm reg_an (a_rm,a_sign,a_exp10,a_is_nan,a_is_inf,a_inf_nan_frac,a_z48,clk,clrn,e, n_rm,n_sign,
    n_exp10,n_is_nan,n_is_inf,n_inf_nan_frac,n_z48);
    // exe3: normalization stage
    fmul_norm mul3 (n_rm,n_sign,n_exp10,n_is_nan,n_is_inf,n_inf_nan_frac,n_z48,s);
endmodule

module fmul_mul (a,b,sign,exp10,s_is_nan,s_is_inf,inf_nan_frac,z_sum,
    z_carry,z8); // mul stage
    input [31:0] a, b;
    output [39:0] z_sum;
    output [39:0] z_carry;
    output [22:0] inf_nan_frac;
    output [9:0] exp10;
    output [7:0] z8;
    output sign;
    output s_is_nan;
    output s_is_inf;
    
    wire a_expo_is_00 = ~|a[30:23]; // exp = 00
    wire b_expo_is_00 = ~|b[30:23];
    wire a_expo_is_ff = &a[30:23]; // exp = ff
    wire b_expo_is_ff = &b[30:23];
    wire a_frac_is_00 = ~|a[22:0]; // frac = 0
    wire b_frac_is_00 = ~|b[22:0];
    wire a_is_inf = a_expo_is_ff & a_frac_is_00;
    wire b_is_inf = b_expo_is_ff & b_frac_is_00;
    wire a_is_nan = a_expo_is_ff & ~a_frac_is_00;
    wire b_is_nan = b_expo_is_ff & ~b_frac_is_00;
    wire a_is_0 = a_expo_is_00 & a_frac_is_00;
    wire b_is_0 = b_expo_is_00 & b_frac_is_00;
    
    assign s_is_inf = a_is_inf | b_is_inf;
    assign s_is_nan = a_is_nan | (a_is_inf & b_is_0) |
            b_is_nan | (b_is_inf & a_is_0);
    wire [22:0] nan_frac = (a[21:0] > b[21:0])?
            {1'b1,a[21:0]} : {1'b1,b[21:0]};
    assign inf_nan_frac = s_is_nan? nan_frac : 23'h0;
    assign sign = a[31] ^ b[31];
    assign exp10 = {2'h0,a[30:23]} + {2'h0,b[30:23]} - 10'h7f +
                a_expo_is_00 + b_expo_is_00; // -126
    wire [23:0] a_frac24 = {~a_expo_is_00,a[22:0]};
    wire [23:0] b_frac24 = {~b_expo_is_00,b[22:0]};
    wallace_24x24 wt24 (a_frac24,b_frac24,z_sum,z_carry,z8);
endmodule

module reg_mul_add (m_rm,m_sign,m_exp10,m_is_nan,m_is_inf,m_inf_nan_frac,
                    m_sum,m_carry,m_z8,clk,clrn,e,a_rm,a_sign,a_exp10,
                    a_is_nan,a_is_inf,a_inf_nan_frac,a_sum,a_carry,a_z8);
    input [39:0] m_sum; // partial mul stage
    input [39:0] m_carry;
    input [22:0] m_inf_nan_frac;
    input [9:0] m_exp10;
    input [7:0] m_z8;
    input [1:0] m_rm;
    input m_sign;
    input m_is_nan;
    input m_is_inf;
    input e; // enable
    input clk, clrn; // clock and reset
    output reg [39:0] a_sum; // addition stage
    output reg [39:0] a_carry;
    output reg [22:0] a_inf_nan_frac;
    output reg [9:0] a_exp10;
    output reg [7:0] a_z8;
    output reg [1:0] a_rm;
    output reg a_sign;
    output reg a_is_nan;
    output reg a_is_inf;
    
    always @ (posedge clk or negedge clrn) begin
        if (!clrn) begin
            a_rm <= 0;
            a_sign <= 0;
            a_exp10 <= 0;
            a_is_nan <= 0;
            a_is_inf <= 0;
            a_inf_nan_frac <= 0;
            a_sum <= 0;
            a_carry <= 0;
            a_z8 <= 0;
        end else if (e) begin
            a_rm <= m_rm;
            a_sign <= m_sign;
            a_exp10 <= m_exp10;
            a_is_nan <= m_is_nan;
            a_is_inf <= m_is_inf;
            a_inf_nan_frac <= m_inf_nan_frac;
            a_sum <= m_sum;
            a_carry <= m_carry;
            a_z8 <= m_z8;
        end
    end
endmodule


module fmul_add (z_sum,z_carry,z); // fmul add
    input [39:0] z_sum;
    input [39:0] z_carry;
    output [47:8] z;
    assign z = z_sum + z_carry;
endmodule

module reg_add_norm (a_rm,a_sign,a_exp10,a_is_nan,a_is_inf,a_inf_nan_frac,
                                a_z48,clk,clrn,e,n_rm,n_sign,n_exp10,n_is_nan,
                                n_is_inf,n_inf_nan_frac,n_z48); // pipeline register
    input [47:0] a_z48; // addition stage
    input [22:0] a_inf_nan_frac;
    input [9:0] a_exp10;
    input [1:0] a_rm;
    input a_sign;
    input a_is_nan;
    input a_is_inf;
    input e; // e: enable
    input clk, clrn; // clock and reset
    output reg [47:0] n_z48; // normalization stage
    output reg [22:0] n_inf_nan_frac;
    output reg [9:0] n_exp10;
    output reg [1:0] n_rm;
    output reg n_sign;
    output reg n_is_nan;
    output reg n_is_inf;

    always @ (posedge clk or negedge clrn) begin
        if (!clrn) begin
            n_rm <= 0;
            n_sign <= 0;
            n_exp10 <= 0;
            n_is_nan <= 0;
            n_is_inf <= 0;
            n_inf_nan_frac <= 0;
            n_z48 <= 0;
        end else if (e) begin
            n_rm <= a_rm;
            n_sign <= a_sign;
            n_exp10 <= a_exp10;
            n_is_nan <= a_is_nan;
            n_is_inf <= a_is_inf;
            n_inf_nan_frac <= a_inf_nan_frac;
            n_z48 <= a_z48;
        end
    end
endmodule


module fmul_norm (rm,sign,exp10,is_nan,is_inf,inf_nan_frac,z,s);// fmul norm
    input [47:0] z; // xx.xxxxxxxxxxxxxxxxxxxxxxxxxx...
    input [22:0] inf_nan_frac;
    input [9:0] exp10;
    input [1:0] rm;
    input sign;
    input is_nan;
    input is_inf;
    output [31:0] s;
    
    wire [46:0] z5,z4,z3,z2,z1,z0; // x.xxxxxxxxxxxxxxxxxxxxxxxxxx...
    wire [5:0] zeros;
    assign zeros[5] = ~|z[46:15]; // 32-bit 0
    assign z5 = zeros[5]? {z[14:0],32'b0} : z[46:0];
    assign zeros[4] = ~|z5[46:31]; // 16-bit 0
    assign z4 = zeros[4]? {z5[30:0],16'b0} : z5;
    assign zeros[3] = ~|z4[46:39]; // 8-bit 0
    assign z3 = zeros[3]? {z4[38:0], 8'b0} : z4;
    assign zeros[2] = ~|z3[46:43]; // 4-bit 0
    assign z2 = zeros[2]? {z3[42:0], 4'b0} : z3;
    assign zeros[1] = ~|z2[46:45]; // 2-bit 0
    assign z1 = zeros[1]? {z2[44:0], 2'b0} : z2;
    assign zeros[0] = ~z1[46]; // 1-bit 0
    assign z0 = zeros[0]? {z1[45:0], 1'b0} : z1;
    reg [46:0] frac0; // temporary fraction
    reg [9:0] exp0; // temporary exponent
    
    always @ * begin
        if (z[47]) begin // 1x.xxxxxxxxxxxxxxxxxxxxxxxx...
            exp0 = exp10 + 10'h1;
            frac0 = z[47:1]; // 1.xxxxxxxxxxxxxxxxxxxxxxxx...
        end else begin
            if (!exp10[9] && (exp10[8:0] > zeros) && z0[46]) begin
                exp0 = exp10 - zeros;
                frac0 = z0; // 1.xxxxxxxxxxxxxxxxxxxxxxxx...
            end else begin // is a denormalized number or 0
                exp0 = 0;
                if (!exp10[9] && (exp10 != 0)) //e>0
                    frac0 = z[46:0] << (exp10 - 10'h1); // e-127 -> -126
                else frac0 = z[46:0] >> (10'h1 - exp10); // e = 0 or neg
            end
        end
    end
    
    wire [26:0] frac = {frac0[46:21],|frac0[20:0]}; // x.xx...xx grs
    wire frac_plus_1 = // for rounding
    ~rm[1] & ~rm[0] & frac0[2] & (frac0[1] | frac0[0]) |
    ~rm[1] & ~rm[0] & frac0[2] & ~frac0[1] & ~frac0[0] & frac0[3] |
    ~rm[1] & rm[0] & (frac0[2] | frac0[1] | frac0[0]) & sign |
    rm[1] & ~rm[0] & (frac0[2] | frac0[1] | frac0[0]) & ~sign;
    wire [24:0] frac_round = {1'b0,frac[26:3]} + frac_plus_1;
    wire [9:0] exp1 = frac_round[24]? exp0 + 10'h1 : exp0;
    wire overflow = (exp0 >= 10'h0ff) | (exp1 >= 10'h0ff);
    
    assign s = final_result(overflow, rm, sign, is_nan, is_inf, exp1[7:0],
                frac_round[22:0], inf_nan_frac);
    
    function [31:0] final_result;
        input overflow;
        input [1:0] rm;
        input sign, is_nan, is_inf;
        input [7:0] exponent;
        input [22:0] fraction,inf_nan_frac;
        
        casex ({overflow,rm,sign,is_nan,is_inf})
            6'b1_00_x_0_x : final_result = {sign,8'hff,23'h000000}; // inf
            6'b1_01_0_0_x : final_result = {sign,8'hfe,23'h7fffff}; // max
            6'b1_01_1_0_x : final_result = {sign,8'hff,23'h000000}; // inf
            6'b1_10_0_0_x : final_result = {sign,8'hff,23'h000000}; // inf
            6'b1_10_1_0_x : final_result = {sign,8'hfe,23'h7fffff}; // max
            6'b1_11_x_0_x : final_result = {sign,8'hfe,23'h7fffff}; // max
            6'b0_xx_x_0_0 : final_result = {sign,exponent,fraction}; // nor
            6'bx_xx_x_1_x : final_result = {1'b1,8'hff,inf_nan_frac}; // nan
            6'bx_xx_x_0_1 : final_result = {sign,8'hff,inf_nan_frac}; // inf
            default : final_result = {sign,8'h00,23'h000000}; // 0
        endcase
    endfunction
endmodule